module FSK_demodulator (
    input wire sys_clk,         // 系统时钟
    input wire rst_n,           // 复位信号 (低电平有效)
    input wire [7:0] phase,     // 当前相位 (0-255)
    input wire signed [7:0] signal, // 输入信号 (显式声明为 signed)
    output reg sign             // 解调输出 (1 或 0)
);

    // 定义中间变量
    reg signed [7:0] sin_val1;
    reg signed [7:0] sin_val2;
    
    // 定义累加器 (24位足够容纳 256 * 8bit * 8bit)
    reg signed [23:0] correlation1;
    reg signed [23:0] correlation2;

    // ============================================================
    // 1. 查找表函数 (ROM 1)
    // ============================================================
    function signed [7:0] get_sin_table1;
        input [7:0] addr;
        begin
            case (addr)
                8'd0: get_sin_table1 = -8'sd1;
                8'd1: get_sin_table1 = 8'sd3;
                8'd2: get_sin_table1 = 8'sd6;
                8'd3: get_sin_table1 = 8'sd9;
                8'd4: get_sin_table1 = 8'sd12;
                8'd5: get_sin_table1 = 8'sd15;
                8'd6: get_sin_table1 = 8'sd18;
                8'd7: get_sin_table1 = 8'sd21;
                8'd8: get_sin_table1 = 8'sd24;
                8'd9: get_sin_table1 = 8'sd28;
                8'd10: get_sin_table1 = 8'sd31;
                8'd11: get_sin_table1 = 8'sd34;
                8'd12: get_sin_table1 = 8'sd37;
                8'd13: get_sin_table1 = 8'sd40;
                8'd14: get_sin_table1 = 8'sd43;
                8'd15: get_sin_table1 = 8'sd46;
                8'd16: get_sin_table1 = 8'sd48;
                8'd17: get_sin_table1 = 8'sd51;
                8'd18: get_sin_table1 = 8'sd54;
                8'd19: get_sin_table1 = 8'sd57;
                8'd20: get_sin_table1 = 8'sd60;
                8'd21: get_sin_table1 = 8'sd63;
                8'd22: get_sin_table1 = 8'sd65;
                8'd23: get_sin_table1 = 8'sd68;
                8'd24: get_sin_table1 = 8'sd71;
                8'd25: get_sin_table1 = 8'sd73;
                8'd26: get_sin_table1 = 8'sd76;
                8'd27: get_sin_table1 = 8'sd78;
                8'd28: get_sin_table1 = 8'sd81;
                8'd29: get_sin_table1 = 8'sd83;
                8'd30: get_sin_table1 = 8'sd85;
                8'd31: get_sin_table1 = 8'sd88;
                8'd32: get_sin_table1 = 8'sd90;
                8'd33: get_sin_table1 = 8'sd92;
                8'd34: get_sin_table1 = 8'sd94;
                8'd35: get_sin_table1 = 8'sd96;
                8'd36: get_sin_table1 = 8'sd98;
                8'd37: get_sin_table1 = 8'sd100;
                8'd38: get_sin_table1 = 8'sd102;
                8'd39: get_sin_table1 = 8'sd104;
                8'd40: get_sin_table1 = 8'sd106;
                8'd41: get_sin_table1 = 8'sd108;
                8'd42: get_sin_table1 = 8'sd109;
                8'd43: get_sin_table1 = 8'sd111;
                8'd44: get_sin_table1 = 8'sd112;
                8'd45: get_sin_table1 = 8'sd114;
                8'd46: get_sin_table1 = 8'sd115;
                8'd47: get_sin_table1 = 8'sd117;
                8'd48: get_sin_table1 = 8'sd118;
                8'd49: get_sin_table1 = 8'sd119;
                8'd50: get_sin_table1 = 8'sd120;
                8'd51: get_sin_table1 = 8'sd121;
                8'd52: get_sin_table1 = 8'sd122;
                8'd53: get_sin_table1 = 8'sd123;
                8'd54: get_sin_table1 = 8'sd124;
                8'd55: get_sin_table1 = 8'sd124;
                8'd56: get_sin_table1 = 8'sd125;
                8'd57: get_sin_table1 = 8'sd126;
                8'd58: get_sin_table1 = 8'sd126;
                8'd59: get_sin_table1 = 8'sd127;
                8'd60: get_sin_table1 = 8'sd127;
                8'd61: get_sin_table1 = 8'sd127;
                8'd62: get_sin_table1 = 8'sd127;
                8'd63: get_sin_table1 = 8'sd127;
                8'd64: get_sin_table1 = 8'sd127;
                8'd65: get_sin_table1 = 8'sd127;
                8'd66: get_sin_table1 = 8'sd127;
                8'd67: get_sin_table1 = 8'sd127;
                8'd68: get_sin_table1 = 8'sd127;
                8'd69: get_sin_table1 = 8'sd127;
                8'd70: get_sin_table1 = 8'sd126;
                8'd71: get_sin_table1 = 8'sd126;
                8'd72: get_sin_table1 = 8'sd125;
                8'd73: get_sin_table1 = 8'sd124;
                8'd74: get_sin_table1 = 8'sd124;
                8'd75: get_sin_table1 = 8'sd123;
                8'd76: get_sin_table1 = 8'sd122;
                8'd77: get_sin_table1 = 8'sd121;
                8'd78: get_sin_table1 = 8'sd120;
                8'd79: get_sin_table1 = 8'sd119;
                8'd80: get_sin_table1 = 8'sd118;
                8'd81: get_sin_table1 = 8'sd117;
                8'd82: get_sin_table1 = 8'sd115;
                8'd83: get_sin_table1 = 8'sd114;
                8'd84: get_sin_table1 = 8'sd112;
                8'd85: get_sin_table1 = 8'sd111;
                8'd86: get_sin_table1 = 8'sd109;
                8'd87: get_sin_table1 = 8'sd108;
                8'd88: get_sin_table1 = 8'sd106;
                8'd89: get_sin_table1 = 8'sd104;
                8'd90: get_sin_table1 = 8'sd102;
                8'd91: get_sin_table1 = 8'sd100;
                8'd92: get_sin_table1 = 8'sd98;
                8'd93: get_sin_table1 = 8'sd96;
                8'd94: get_sin_table1 = 8'sd94;
                8'd95: get_sin_table1 = 8'sd92;
                8'd96: get_sin_table1 = 8'sd90;
                8'd97: get_sin_table1 = 8'sd88;
                8'd98: get_sin_table1 = 8'sd85;
                8'd99: get_sin_table1 = 8'sd83;
                8'd100: get_sin_table1 = 8'sd81;
                8'd101: get_sin_table1 = 8'sd78;
                8'd102: get_sin_table1 = 8'sd76;
                8'd103: get_sin_table1 = 8'sd73;
                8'd104: get_sin_table1 = 8'sd71;
                8'd105: get_sin_table1 = 8'sd68;
                8'd106: get_sin_table1 = 8'sd65;
                8'd107: get_sin_table1 = 8'sd63;
                8'd108: get_sin_table1 = 8'sd60;
                8'd109: get_sin_table1 = 8'sd57;
                8'd110: get_sin_table1 = 8'sd54;
                8'd111: get_sin_table1 = 8'sd51;
                8'd112: get_sin_table1 = 8'sd48;
                8'd113: get_sin_table1 = 8'sd46;
                8'd114: get_sin_table1 = 8'sd43;
                8'd115: get_sin_table1 = 8'sd40;
                8'd116: get_sin_table1 = 8'sd37;
                8'd117: get_sin_table1 = 8'sd34;
                8'd118: get_sin_table1 = 8'sd31;
                8'd119: get_sin_table1 = 8'sd28;
                8'd120: get_sin_table1 = 8'sd24;
                8'd121: get_sin_table1 = 8'sd21;
                8'd122: get_sin_table1 = 8'sd18;
                8'd123: get_sin_table1 = 8'sd15;
                8'd124: get_sin_table1 = 8'sd12;
                8'd125: get_sin_table1 = 8'sd9;
                8'd126: get_sin_table1 = 8'sd6;
                8'd127: get_sin_table1 = 8'sd3;
                8'd128: get_sin_table1 = 8'sd0;
                8'd129: get_sin_table1 = -8'sd4;
                8'd130: get_sin_table1 = -8'sd7;
                8'd131: get_sin_table1 = -8'sd10;
                8'd132: get_sin_table1 = -8'sd13;
                8'd133: get_sin_table1 = -8'sd16;
                8'd134: get_sin_table1 = -8'sd19;
                8'd135: get_sin_table1 = -8'sd22;
                8'd136: get_sin_table1 = -8'sd25;
                8'd137: get_sin_table1 = -8'sd29;
                8'd138: get_sin_table1 = -8'sd32;
                8'd139: get_sin_table1 = -8'sd35;
                8'd140: get_sin_table1 = -8'sd38;
                8'd141: get_sin_table1 = -8'sd41;
                8'd142: get_sin_table1 = -8'sd44;
                8'd143: get_sin_table1 = -8'sd47;
                8'd144: get_sin_table1 = -8'sd49;
                8'd145: get_sin_table1 = -8'sd52;
                8'd146: get_sin_table1 = -8'sd55;
                8'd147: get_sin_table1 = -8'sd58;
                8'd148: get_sin_table1 = -8'sd61;
                8'd149: get_sin_table1 = -8'sd64;
                8'd150: get_sin_table1 = -8'sd66;
                8'd151: get_sin_table1 = -8'sd69;
                8'd152: get_sin_table1 = -8'sd72;
                8'd153: get_sin_table1 = -8'sd74;
                8'd154: get_sin_table1 = -8'sd77;
                8'd155: get_sin_table1 = -8'sd79;
                8'd156: get_sin_table1 = -8'sd82;
                8'd157: get_sin_table1 = -8'sd84;
                8'd158: get_sin_table1 = -8'sd86;
                8'd159: get_sin_table1 = -8'sd89;
                8'd160: get_sin_table1 = -8'sd91;
                8'd161: get_sin_table1 = -8'sd93;
                8'd162: get_sin_table1 = -8'sd95;
                8'd163: get_sin_table1 = -8'sd97;
                8'd164: get_sin_table1 = -8'sd99;
                8'd165: get_sin_table1 = -8'sd101;
                8'd166: get_sin_table1 = -8'sd103;
                8'd167: get_sin_table1 = -8'sd105;
                8'd168: get_sin_table1 = -8'sd107;
                8'd169: get_sin_table1 = -8'sd109;
                8'd170: get_sin_table1 = -8'sd110;
                8'd171: get_sin_table1 = -8'sd112;
                8'd172: get_sin_table1 = -8'sd113;
                8'd173: get_sin_table1 = -8'sd115;
                8'd174: get_sin_table1 = -8'sd116;
                8'd175: get_sin_table1 = -8'sd118;
                8'd176: get_sin_table1 = -8'sd119;
                8'd177: get_sin_table1 = -8'sd120;
                8'd178: get_sin_table1 = -8'sd121;
                8'd179: get_sin_table1 = -8'sd122;
                8'd180: get_sin_table1 = -8'sd123;
                8'd181: get_sin_table1 = -8'sd124;
                8'd182: get_sin_table1 = -8'sd125;
                8'd183: get_sin_table1 = -8'sd125;
                8'd184: get_sin_table1 = -8'sd126;
                8'd185: get_sin_table1 = -8'sd127;
                8'd186: get_sin_table1 = -8'sd127;
                8'd187: get_sin_table1 = -8'sd128;
                8'd188: get_sin_table1 = -8'sd128;
                8'd189: get_sin_table1 = -8'sd128;
                8'd190: get_sin_table1 = -8'sd128;
                8'd191: get_sin_table1 = -8'sd128;
                8'd192: get_sin_table1 = -8'sd129;
                8'd193: get_sin_table1 = -8'sd128;
                8'd194: get_sin_table1 = -8'sd128;
                8'd195: get_sin_table1 = -8'sd128;
                8'd196: get_sin_table1 = -8'sd128;
                8'd197: get_sin_table1 = -8'sd128;
                8'd198: get_sin_table1 = -8'sd127;
                8'd199: get_sin_table1 = -8'sd127;
                8'd200: get_sin_table1 = -8'sd126;
                8'd201: get_sin_table1 = -8'sd125;
                8'd202: get_sin_table1 = -8'sd125;
                8'd203: get_sin_table1 = -8'sd124;
                8'd204: get_sin_table1 = -8'sd123;
                8'd205: get_sin_table1 = -8'sd122;
                8'd206: get_sin_table1 = -8'sd121;
                8'd207: get_sin_table1 = -8'sd120;
                8'd208: get_sin_table1 = -8'sd119;
                8'd209: get_sin_table1 = -8'sd118;
                8'd210: get_sin_table1 = -8'sd116;
                8'd211: get_sin_table1 = -8'sd115;
                8'd212: get_sin_table1 = -8'sd113;
                8'd213: get_sin_table1 = -8'sd112;
                8'd214: get_sin_table1 = -8'sd110;
                8'd215: get_sin_table1 = -8'sd109;
                8'd216: get_sin_table1 = -8'sd107;
                8'd217: get_sin_table1 = -8'sd105;
                8'd218: get_sin_table1 = -8'sd103;
                8'd219: get_sin_table1 = -8'sd101;
                8'd220: get_sin_table1 = -8'sd99;
                8'd221: get_sin_table1 = -8'sd97;
                8'd222: get_sin_table1 = -8'sd95;
                8'd223: get_sin_table1 = -8'sd93;
                8'd224: get_sin_table1 = -8'sd91;
                8'd225: get_sin_table1 = -8'sd89;
                8'd226: get_sin_table1 = -8'sd86;
                8'd227: get_sin_table1 = -8'sd84;
                8'd228: get_sin_table1 = -8'sd82;
                8'd229: get_sin_table1 = -8'sd79;
                8'd230: get_sin_table1 = -8'sd77;
                8'd231: get_sin_table1 = -8'sd74;
                8'd232: get_sin_table1 = -8'sd72;
                8'd233: get_sin_table1 = -8'sd69;
                8'd234: get_sin_table1 = -8'sd66;
                8'd235: get_sin_table1 = -8'sd64;
                8'd236: get_sin_table1 = -8'sd61;
                8'd237: get_sin_table1 = -8'sd58;
                8'd238: get_sin_table1 = -8'sd55;
                8'd239: get_sin_table1 = -8'sd52;
                8'd240: get_sin_table1 = -8'sd49;
                8'd241: get_sin_table1 = -8'sd47;
                8'd242: get_sin_table1 = -8'sd44;
                8'd243: get_sin_table1 = -8'sd41;
                8'd244: get_sin_table1 = -8'sd38;
                8'd245: get_sin_table1 = -8'sd35;
                8'd246: get_sin_table1 = -8'sd32;
                8'd247: get_sin_table1 = -8'sd29;
                8'd248: get_sin_table1 = -8'sd25;
                8'd249: get_sin_table1 = -8'sd22;
                8'd250: get_sin_table1 = -8'sd19;
                8'd251: get_sin_table1 = -8'sd16;
                8'd252: get_sin_table1 = -8'sd13;
                8'd253: get_sin_table1 = -8'sd10;
                8'd254: get_sin_table1 = -8'sd7;
                8'd255: get_sin_table1 = -8'sd4;
                default: get_sin_table1 = 8'sd0;
            endcase
        end
    endfunction

    // ============================================================
    // 2. 查找表函数 (ROM 2)
    // ============================================================
    function signed [7:0] get_sin_table2;
        input [7:0] addr;
        begin
            case (addr)
                8'd0: get_sin_table2 = -8'sd1;
                8'd1: get_sin_table2 = 8'sd6;
                8'd2: get_sin_table2 = 8'sd12;
                8'd3: get_sin_table2 = 8'sd18;
                8'd4: get_sin_table2 = 8'sd24;
                8'd5: get_sin_table2 = 8'sd31;
                8'd6: get_sin_table2 = 8'sd37;
                8'd7: get_sin_table2 = 8'sd43;
                8'd8: get_sin_table2 = 8'sd48;
                8'd9: get_sin_table2 = 8'sd54;
                8'd10: get_sin_table2 = 8'sd60;
                8'd11: get_sin_table2 = 8'sd65;
                8'd12: get_sin_table2 = 8'sd71;
                8'd13: get_sin_table2 = 8'sd76;
                8'd14: get_sin_table2 = 8'sd81;
                8'd15: get_sin_table2 = 8'sd85;
                8'd16: get_sin_table2 = 8'sd90;
                8'd17: get_sin_table2 = 8'sd94;
                8'd18: get_sin_table2 = 8'sd98;
                8'd19: get_sin_table2 = 8'sd102;
                8'd20: get_sin_table2 = 8'sd106;
                8'd21: get_sin_table2 = 8'sd109;
                8'd22: get_sin_table2 = 8'sd112;
                8'd23: get_sin_table2 = 8'sd115;
                8'd24: get_sin_table2 = 8'sd118;
                8'd25: get_sin_table2 = 8'sd120;
                8'd26: get_sin_table2 = 8'sd122;
                8'd27: get_sin_table2 = 8'sd124;
                8'd28: get_sin_table2 = 8'sd125;
                8'd29: get_sin_table2 = 8'sd126;
                8'd30: get_sin_table2 = 8'sd127;
                8'd31: get_sin_table2 = 8'sd127;
                8'd32: get_sin_table2 = 8'sd127;
                8'd33: get_sin_table2 = 8'sd127;
                8'd34: get_sin_table2 = 8'sd127;
                8'd35: get_sin_table2 = 8'sd126;
                8'd36: get_sin_table2 = 8'sd125;
                8'd37: get_sin_table2 = 8'sd124;
                8'd38: get_sin_table2 = 8'sd122;
                8'd39: get_sin_table2 = 8'sd120;
                8'd40: get_sin_table2 = 8'sd118;
                8'd41: get_sin_table2 = 8'sd115;
                8'd42: get_sin_table2 = 8'sd112;
                8'd43: get_sin_table2 = 8'sd109;
                8'd44: get_sin_table2 = 8'sd106;
                8'd45: get_sin_table2 = 8'sd102;
                8'd46: get_sin_table2 = 8'sd98;
                8'd47: get_sin_table2 = 8'sd94;
                8'd48: get_sin_table2 = 8'sd90;
                8'd49: get_sin_table2 = 8'sd85;
                8'd50: get_sin_table2 = 8'sd81;
                8'd51: get_sin_table2 = 8'sd76;
                8'd52: get_sin_table2 = 8'sd71;
                8'd53: get_sin_table2 = 8'sd65;
                8'd54: get_sin_table2 = 8'sd60;
                8'd55: get_sin_table2 = 8'sd54;
                8'd56: get_sin_table2 = 8'sd48;
                8'd57: get_sin_table2 = 8'sd43;
                8'd58: get_sin_table2 = 8'sd37;
                8'd59: get_sin_table2 = 8'sd31;
                8'd60: get_sin_table2 = 8'sd24;
                8'd61: get_sin_table2 = 8'sd18;
                8'd62: get_sin_table2 = 8'sd12;
                8'd63: get_sin_table2 = 8'sd6;
                8'd64: get_sin_table2 = 8'sd0;
                8'd65: get_sin_table2 = -8'sd7;
                8'd66: get_sin_table2 = -8'sd13;
                8'd67: get_sin_table2 = -8'sd19;
                8'd68: get_sin_table2 = -8'sd25;
                8'd69: get_sin_table2 = -8'sd32;
                8'd70: get_sin_table2 = -8'sd38;
                8'd71: get_sin_table2 = -8'sd44;
                8'd72: get_sin_table2 = -8'sd49;
                8'd73: get_sin_table2 = -8'sd55;
                8'd74: get_sin_table2 = -8'sd61;
                8'd75: get_sin_table2 = -8'sd66;
                8'd76: get_sin_table2 = -8'sd72;
                8'd77: get_sin_table2 = -8'sd77;
                8'd78: get_sin_table2 = -8'sd82;
                8'd79: get_sin_table2 = -8'sd86;
                8'd80: get_sin_table2 = -8'sd91;
                8'd81: get_sin_table2 = -8'sd95;
                8'd82: get_sin_table2 = -8'sd99;
                8'd83: get_sin_table2 = -8'sd103;
                8'd84: get_sin_table2 = -8'sd107;
                8'd85: get_sin_table2 = -8'sd110;
                8'd86: get_sin_table2 = -8'sd113;
                8'd87: get_sin_table2 = -8'sd116;
                8'd88: get_sin_table2 = -8'sd119;
                8'd89: get_sin_table2 = -8'sd121;
                8'd90: get_sin_table2 = -8'sd123;
                8'd91: get_sin_table2 = -8'sd125;
                8'd92: get_sin_table2 = -8'sd126;
                8'd93: get_sin_table2 = -8'sd127;
                8'd94: get_sin_table2 = -8'sd128;
                8'd95: get_sin_table2 = -8'sd128;
                8'd96: get_sin_table2 = -8'sd129;
                8'd97: get_sin_table2 = -8'sd128;
                8'd98: get_sin_table2 = -8'sd128;
                8'd99: get_sin_table2 = -8'sd127;
                8'd100: get_sin_table2 = -8'sd126;
                8'd101: get_sin_table2 = -8'sd125;
                8'd102: get_sin_table2 = -8'sd123;
                8'd103: get_sin_table2 = -8'sd121;
                8'd104: get_sin_table2 = -8'sd119;
                8'd105: get_sin_table2 = -8'sd116;
                8'd106: get_sin_table2 = -8'sd113;
                8'd107: get_sin_table2 = -8'sd110;
                8'd108: get_sin_table2 = -8'sd107;
                8'd109: get_sin_table2 = -8'sd103;
                8'd110: get_sin_table2 = -8'sd99;
                8'd111: get_sin_table2 = -8'sd95;
                8'd112: get_sin_table2 = -8'sd91;
                8'd113: get_sin_table2 = -8'sd86;
                8'd114: get_sin_table2 = -8'sd82;
                8'd115: get_sin_table2 = -8'sd77;
                8'd116: get_sin_table2 = -8'sd72;
                8'd117: get_sin_table2 = -8'sd66;
                8'd118: get_sin_table2 = -8'sd61;
                8'd119: get_sin_table2 = -8'sd55;
                8'd120: get_sin_table2 = -8'sd49;
                8'd121: get_sin_table2 = -8'sd44;
                8'd122: get_sin_table2 = -8'sd38;
                8'd123: get_sin_table2 = -8'sd32;
                8'd124: get_sin_table2 = -8'sd25;
                8'd125: get_sin_table2 = -8'sd19;
                8'd126: get_sin_table2 = -8'sd13;
                8'd127: get_sin_table2 = -8'sd7;
                8'd128: get_sin_table2 = -8'sd1;
                8'd129: get_sin_table2 = 8'sd6;
                8'd130: get_sin_table2 = 8'sd12;
                8'd131: get_sin_table2 = 8'sd18;
                8'd132: get_sin_table2 = 8'sd24;
                8'd133: get_sin_table2 = 8'sd31;
                8'd134: get_sin_table2 = 8'sd37;
                8'd135: get_sin_table2 = 8'sd43;
                8'd136: get_sin_table2 = 8'sd48;
                8'd137: get_sin_table2 = 8'sd54;
                8'd138: get_sin_table2 = 8'sd60;
                8'd139: get_sin_table2 = 8'sd65;
                8'd140: get_sin_table2 = 8'sd71;
                8'd141: get_sin_table2 = 8'sd76;
                8'd142: get_sin_table2 = 8'sd81;
                8'd143: get_sin_table2 = 8'sd85;
                8'd144: get_sin_table2 = 8'sd90;
                8'd145: get_sin_table2 = 8'sd94;
                8'd146: get_sin_table2 = 8'sd98;
                8'd147: get_sin_table2 = 8'sd102;
                8'd148: get_sin_table2 = 8'sd106;
                8'd149: get_sin_table2 = 8'sd109;
                8'd150: get_sin_table2 = 8'sd112;
                8'd151: get_sin_table2 = 8'sd115;
                8'd152: get_sin_table2 = 8'sd118;
                8'd153: get_sin_table2 = 8'sd120;
                8'd154: get_sin_table2 = 8'sd122;
                8'd155: get_sin_table2 = 8'sd124;
                8'd156: get_sin_table2 = 8'sd125;
                8'd157: get_sin_table2 = 8'sd126;
                8'd158: get_sin_table2 = 8'sd127;
                8'd159: get_sin_table2 = 8'sd127;
                8'd160: get_sin_table2 = 8'sd127;
                8'd161: get_sin_table2 = 8'sd127;
                8'd162: get_sin_table2 = 8'sd127;
                8'd163: get_sin_table2 = 8'sd126;
                8'd164: get_sin_table2 = 8'sd125;
                8'd165: get_sin_table2 = 8'sd124;
                8'd166: get_sin_table2 = 8'sd122;
                8'd167: get_sin_table2 = 8'sd120;
                8'd168: get_sin_table2 = 8'sd118;
                8'd169: get_sin_table2 = 8'sd115;
                8'd170: get_sin_table2 = 8'sd112;
                8'd171: get_sin_table2 = 8'sd109;
                8'd172: get_sin_table2 = 8'sd106;
                8'd173: get_sin_table2 = 8'sd102;
                8'd174: get_sin_table2 = 8'sd98;
                8'd175: get_sin_table2 = 8'sd94;
                8'd176: get_sin_table2 = 8'sd90;
                8'd177: get_sin_table2 = 8'sd85;
                8'd178: get_sin_table2 = 8'sd81;
                8'd179: get_sin_table2 = 8'sd76;
                8'd180: get_sin_table2 = 8'sd71;
                8'd181: get_sin_table2 = 8'sd65;
                8'd182: get_sin_table2 = 8'sd60;
                8'd183: get_sin_table2 = 8'sd54;
                8'd184: get_sin_table2 = 8'sd48;
                8'd185: get_sin_table2 = 8'sd43;
                8'd186: get_sin_table2 = 8'sd37;
                8'd187: get_sin_table2 = 8'sd31;
                8'd188: get_sin_table2 = 8'sd24;
                8'd189: get_sin_table2 = 8'sd18;
                8'd190: get_sin_table2 = 8'sd12;
                8'd191: get_sin_table2 = 8'sd6;
                8'd192: get_sin_table2 = 8'sd0;
                8'd193: get_sin_table2 = -8'sd7;
                8'd194: get_sin_table2 = -8'sd13;
                8'd195: get_sin_table2 = -8'sd19;
                8'd196: get_sin_table2 = -8'sd25;
                8'd197: get_sin_table2 = -8'sd32;
                8'd198: get_sin_table2 = -8'sd38;
                8'd199: get_sin_table2 = -8'sd44;
                8'd200: get_sin_table2 = -8'sd49;
                8'd201: get_sin_table2 = -8'sd55;
                8'd202: get_sin_table2 = -8'sd61;
                8'd203: get_sin_table2 = -8'sd66;
                8'd204: get_sin_table2 = -8'sd72;
                8'd205: get_sin_table2 = -8'sd77;
                8'd206: get_sin_table2 = -8'sd82;
                8'd207: get_sin_table2 = -8'sd86;
                8'd208: get_sin_table2 = -8'sd91;
                8'd209: get_sin_table2 = -8'sd95;
                8'd210: get_sin_table2 = -8'sd99;
                8'd211: get_sin_table2 = -8'sd103;
                8'd212: get_sin_table2 = -8'sd107;
                8'd213: get_sin_table2 = -8'sd110;
                8'd214: get_sin_table2 = -8'sd113;
                8'd215: get_sin_table2 = -8'sd116;
                8'd216: get_sin_table2 = -8'sd119;
                8'd217: get_sin_table2 = -8'sd121;
                8'd218: get_sin_table2 = -8'sd123;
                8'd219: get_sin_table2 = -8'sd125;
                8'd220: get_sin_table2 = -8'sd126;
                8'd221: get_sin_table2 = -8'sd127;
                8'd222: get_sin_table2 = -8'sd128;
                8'd223: get_sin_table2 = -8'sd128;
                8'd224: get_sin_table2 = -8'sd129;
                8'd225: get_sin_table2 = -8'sd128;
                8'd226: get_sin_table2 = -8'sd128;
                8'd227: get_sin_table2 = -8'sd127;
                8'd228: get_sin_table2 = -8'sd126;
                8'd229: get_sin_table2 = -8'sd125;
                8'd230: get_sin_table2 = -8'sd123;
                8'd231: get_sin_table2 = -8'sd121;
                8'd232: get_sin_table2 = -8'sd119;
                8'd233: get_sin_table2 = -8'sd116;
                8'd234: get_sin_table2 = -8'sd113;
                8'd235: get_sin_table2 = -8'sd110;
                8'd236: get_sin_table2 = -8'sd107;
                8'd237: get_sin_table2 = -8'sd103;
                8'd238: get_sin_table2 = -8'sd99;
                8'd239: get_sin_table2 = -8'sd95;
                8'd240: get_sin_table2 = -8'sd91;
                8'd241: get_sin_table2 = -8'sd86;
                8'd242: get_sin_table2 = -8'sd82;
                8'd243: get_sin_table2 = -8'sd77;
                8'd244: get_sin_table2 = -8'sd72;
                8'd245: get_sin_table2 = -8'sd66;
                8'd246: get_sin_table2 = -8'sd61;
                8'd247: get_sin_table2 = -8'sd55;
                8'd248: get_sin_table2 = -8'sd49;
                8'd249: get_sin_table2 = -8'sd44;
                8'd250: get_sin_table2 = -8'sd38;
                8'd251: get_sin_table2 = -8'sd32;
                8'd252: get_sin_table2 = -8'sd25;
                8'd253: get_sin_table2 = -8'sd19;
                8'd254: get_sin_table2 = -8'sd13;
                8'd255: get_sin_table2 = -8'sd7;
                default: get_sin_table2 = 8'sd0;
            endcase
        end
    endfunction


    // ============================================================
    // 3. 主逻辑 (完全同步设计)
    // ============================================================
    always @(posedge sys_clk or negedge rst_n) begin
        if (!rst_n) begin
            correlation1 <= 0;
            correlation2 <= 0;
            sign <= 0;
            sin_val1 <= 0;
            sin_val2 <= 0;
        end
        else begin

            sin_val1 <= get_sin_table1(phase);
            sin_val2 <= get_sin_table2(phase);
            
            if (phase == 255) begin

                if (correlation1 > correlation2)
                    sign <= 1;
                else
                    sign <= 0;
            
                correlation1 <= sin_val1 * signal; 
                correlation2 <= sin_val2 * signal;
            end 
            else begin
                // 正常的乘累加运算
                correlation1 <= correlation1 + (sin_val1 * signal);
                correlation2 <= correlation2 + (sin_val2 * signal);
            end
        end
    end

endmodule