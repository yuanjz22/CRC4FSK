module FSK_demodulator (
   input wire clk_sign,
   input wire [7:0] phase,
   input wire [7:0] signal,
   output reg sign
);

   reg signed [7:0] sin_table1 [0:255];
   reg signed [7:0] sin_table2 [0:255];
   reg signed [23:0] correlation1;
   reg signed [23:0] correlation2;

   initial begin
       sin_table1[0] = -1;
       sin_table1[1] = 3;
       sin_table1[2] = 6;
       sin_table1[3] = 9;
       sin_table1[4] = 12;
       sin_table1[5] = 15;
       sin_table1[6] = 18;
       sin_table1[7] = 21;
       sin_table1[8] = 24;
       sin_table1[9] = 28;
       sin_table1[10] = 31;
       sin_table1[11] = 34;
       sin_table1[12] = 37;
       sin_table1[13] = 40;
       sin_table1[14] = 43;
       sin_table1[15] = 46;
       sin_table1[16] = 48;
       sin_table1[17] = 51;
       sin_table1[18] = 54;
       sin_table1[19] = 57;
       sin_table1[20] = 60;
       sin_table1[21] = 63;
       sin_table1[22] = 65;
       sin_table1[23] = 68;
       sin_table1[24] = 71;
       sin_table1[25] = 73;
       sin_table1[26] = 76;
       sin_table1[27] = 78;
       sin_table1[28] = 81;
       sin_table1[29] = 83;
       sin_table1[30] = 85;
       sin_table1[31] = 88;
       sin_table1[32] = 90;
       sin_table1[33] = 92;
       sin_table1[34] = 94;
       sin_table1[35] = 96;
       sin_table1[36] = 98;
       sin_table1[37] = 100;
       sin_table1[38] = 102;
       sin_table1[39] = 104;
       sin_table1[40] = 106;
       sin_table1[41] = 108;
       sin_table1[42] = 109;
       sin_table1[43] = 111;
       sin_table1[44] = 112;
       sin_table1[45] = 114;
       sin_table1[46] = 115;
       sin_table1[47] = 117;
       sin_table1[48] = 118;
       sin_table1[49] = 119;
       sin_table1[50] = 120;
       sin_table1[51] = 121;
       sin_table1[52] = 122;
       sin_table1[53] = 123;
       sin_table1[54] = 124;
       sin_table1[55] = 124;
       sin_table1[56] = 125;
       sin_table1[57] = 126;
       sin_table1[58] = 126;
       sin_table1[59] = 127;
       sin_table1[60] = 127;
       sin_table1[61] = 127;
       sin_table1[62] = 127;
       sin_table1[63] = 127;
       sin_table1[64] = 127;
       sin_table1[65] = 127;
       sin_table1[66] = 127;
       sin_table1[67] = 127;
       sin_table1[68] = 127;
       sin_table1[69] = 127;
       sin_table1[70] = 126;
       sin_table1[71] = 126;
       sin_table1[72] = 125;
       sin_table1[73] = 124;
       sin_table1[74] = 124;
       sin_table1[75] = 123;
       sin_table1[76] = 122;
       sin_table1[77] = 121;
       sin_table1[78] = 120;
       sin_table1[79] = 119;
       sin_table1[80] = 118;
       sin_table1[81] = 117;
       sin_table1[82] = 115;
       sin_table1[83] = 114;
       sin_table1[84] = 112;
       sin_table1[85] = 111;
       sin_table1[86] = 109;
       sin_table1[87] = 108;
       sin_table1[88] = 106;
       sin_table1[89] = 104;
       sin_table1[90] = 102;
       sin_table1[91] = 100;
       sin_table1[92] = 98;
       sin_table1[93] = 96;
       sin_table1[94] = 94;
       sin_table1[95] = 92;
       sin_table1[96] = 90;
       sin_table1[97] = 88;
       sin_table1[98] = 85;
       sin_table1[99] = 83;
       sin_table1[100] = 81;
       sin_table1[101] = 78;
       sin_table1[102] = 76;
       sin_table1[103] = 73;
       sin_table1[104] = 71;
       sin_table1[105] = 68;
       sin_table1[106] = 65;
       sin_table1[107] = 63;
       sin_table1[108] = 60;
       sin_table1[109] = 57;
       sin_table1[110] = 54;
       sin_table1[111] = 51;
       sin_table1[112] = 48;
       sin_table1[113] = 46;
       sin_table1[114] = 43;
       sin_table1[115] = 40;
       sin_table1[116] = 37;
       sin_table1[117] = 34;
       sin_table1[118] = 31;
       sin_table1[119] = 28;
       sin_table1[120] = 24;
       sin_table1[121] = 21;
       sin_table1[122] = 18;
       sin_table1[123] = 15;
       sin_table1[124] = 12;
       sin_table1[125] = 9;
       sin_table1[126] = 6;
       sin_table1[127] = 3;
       sin_table1[128] = 0;
       sin_table1[129] = -4;
       sin_table1[130] = -7;
       sin_table1[131] = -10;
       sin_table1[132] = -13;
       sin_table1[133] = -16;
       sin_table1[134] = -19;
       sin_table1[135] = -22;
       sin_table1[136] = -25;
       sin_table1[137] = -29;
       sin_table1[138] = -32;
       sin_table1[139] = -35;
       sin_table1[140] = -38;
       sin_table1[141] = -41;
       sin_table1[142] = -44;
       sin_table1[143] = -47;
       sin_table1[144] = -49;
       sin_table1[145] = -52;
       sin_table1[146] = -55;
       sin_table1[147] = -58;
       sin_table1[148] = -61;
       sin_table1[149] = -64;
       sin_table1[150] = -66;
       sin_table1[151] = -69;
       sin_table1[152] = -72;
       sin_table1[153] = -74;
       sin_table1[154] = -77;
       sin_table1[155] = -79;
       sin_table1[156] = -82;
       sin_table1[157] = -84;
       sin_table1[158] = -86;
       sin_table1[159] = -89;
       sin_table1[160] = -91;
       sin_table1[161] = -93;
       sin_table1[162] = -95;
       sin_table1[163] = -97;
       sin_table1[164] = -99;
       sin_table1[165] = -101;
       sin_table1[166] = -103;
       sin_table1[167] = -105;
       sin_table1[168] = -107;
       sin_table1[169] = -109;
       sin_table1[170] = -110;
       sin_table1[171] = -112;
       sin_table1[172] = -113;
       sin_table1[173] = -115;
       sin_table1[174] = -116;
       sin_table1[175] = -118;
       sin_table1[176] = -119;
       sin_table1[177] = -120;
       sin_table1[178] = -121;
       sin_table1[179] = -122;
       sin_table1[180] = -123;
       sin_table1[181] = -124;
       sin_table1[182] = -125;
       sin_table1[183] = -125;
       sin_table1[184] = -126;
       sin_table1[185] = -127;
       sin_table1[186] = -127;
       sin_table1[187] = -128;
       sin_table1[188] = -128;
       sin_table1[189] = -128;
       sin_table1[190] = -128;
       sin_table1[191] = -128;
       sin_table1[192] = -129;
       sin_table1[193] = -128;
       sin_table1[194] = -128;
       sin_table1[195] = -128;
       sin_table1[196] = -128;
       sin_table1[197] = -128;
       sin_table1[198] = -127;
       sin_table1[199] = -127;
       sin_table1[200] = -126;
       sin_table1[201] = -125;
       sin_table1[202] = -125;
       sin_table1[203] = -124;
       sin_table1[204] = -123;
       sin_table1[205] = -122;
       sin_table1[206] = -121;
       sin_table1[207] = -120;
       sin_table1[208] = -119;
       sin_table1[209] = -118;
       sin_table1[210] = -116;
       sin_table1[211] = -115;
       sin_table1[212] = -113;
       sin_table1[213] = -112;
       sin_table1[214] = -110;
       sin_table1[215] = -109;
       sin_table1[216] = -107;
       sin_table1[217] = -105;
       sin_table1[218] = -103;
       sin_table1[219] = -101;
       sin_table1[220] = -99;
       sin_table1[221] = -97;
       sin_table1[222] = -95;
       sin_table1[223] = -93;
       sin_table1[224] = -91;
       sin_table1[225] = -89;
       sin_table1[226] = -86;
       sin_table1[227] = -84;
       sin_table1[228] = -82;
       sin_table1[229] = -79;
       sin_table1[230] = -77;
       sin_table1[231] = -74;
       sin_table1[232] = -72;
       sin_table1[233] = -69;
       sin_table1[234] = -66;
       sin_table1[235] = -64;
       sin_table1[236] = -61;
       sin_table1[237] = -58;
       sin_table1[238] = -55;
       sin_table1[239] = -52;
       sin_table1[240] = -49;
       sin_table1[241] = -47;
       sin_table1[242] = -44;
       sin_table1[243] = -41;
       sin_table1[244] = -38;
       sin_table1[245] = -35;
       sin_table1[246] = -32;
       sin_table1[247] = -29;
       sin_table1[248] = -25;
       sin_table1[249] = -22;
       sin_table1[250] = -19;
       sin_table1[251] = -16;
       sin_table1[252] = -13;
       sin_table1[253] = -10;
       sin_table1[254] = -7;
       sin_table1[255] = -4;

       sin_table2[0] = -1;
       sin_table2[1] = 6;
       sin_table2[2] = 12;
       sin_table2[3] = 18;
       sin_table2[4] = 24;
       sin_table2[5] = 31;
       sin_table2[6] = 37;
       sin_table2[7] = 43;
       sin_table2[8] = 48;
       sin_table2[9] = 54;
       sin_table2[10] = 60;
       sin_table2[11] = 65;
       sin_table2[12] = 71;
       sin_table2[13] = 76;
       sin_table2[14] = 81;
       sin_table2[15] = 85;
       sin_table2[16] = 90;
       sin_table2[17] = 94;
       sin_table2[18] = 98;
       sin_table2[19] = 102;
       sin_table2[20] = 106;
       sin_table2[21] = 109;
       sin_table2[22] = 112;
       sin_table2[23] = 115;
       sin_table2[24] = 118;
       sin_table2[25] = 120;
       sin_table2[26] = 122;
       sin_table2[27] = 124;
       sin_table2[28] = 125;
       sin_table2[29] = 126;
       sin_table2[30] = 127;
       sin_table2[31] = 127;
       sin_table2[32] = 127;
       sin_table2[33] = 127;
       sin_table2[34] = 127;
       sin_table2[35] = 126;
       sin_table2[36] = 125;
       sin_table2[37] = 124;
       sin_table2[38] = 122;
       sin_table2[39] = 120;
       sin_table2[40] = 118;
       sin_table2[41] = 115;
       sin_table2[42] = 112;
       sin_table2[43] = 109;
       sin_table2[44] = 106;
       sin_table2[45] = 102;
       sin_table2[46] = 98;
       sin_table2[47] = 94;
       sin_table2[48] = 90;
       sin_table2[49] = 85;
       sin_table2[50] = 81;
       sin_table2[51] = 76;
       sin_table2[52] = 71;
       sin_table2[53] = 65;
       sin_table2[54] = 60;
       sin_table2[55] = 54;
       sin_table2[56] = 48;
       sin_table2[57] = 43;
       sin_table2[58] = 37;
       sin_table2[59] = 31;
       sin_table2[60] = 24;
       sin_table2[61] = 18;
       sin_table2[62] = 12;
       sin_table2[63] = 6;
       sin_table2[64] = 0;
       sin_table2[65] = -7;
       sin_table2[66] = -13;
       sin_table2[67] = -19;
       sin_table2[68] = -25;
       sin_table2[69] = -32;
       sin_table2[70] = -38;
       sin_table2[71] = -44;
       sin_table2[72] = -49;
       sin_table2[73] = -55;
       sin_table2[74] = -61;
       sin_table2[75] = -66;
       sin_table2[76] = -72;
       sin_table2[77] = -77;
       sin_table2[78] = -82;
       sin_table2[79] = -86;
       sin_table2[80] = -91;
       sin_table2[81] = -95;
       sin_table2[82] = -99;
       sin_table2[83] = -103;
       sin_table2[84] = -107;
       sin_table2[85] = -110;
       sin_table2[86] = -113;
       sin_table2[87] = -116;
       sin_table2[88] = -119;
       sin_table2[89] = -121;
       sin_table2[90] = -123;
       sin_table2[91] = -125;
       sin_table2[92] = -126;
       sin_table2[93] = -127;
       sin_table2[94] = -128;
       sin_table2[95] = -128;
       sin_table2[96] = -129;
       sin_table2[97] = -128;
       sin_table2[98] = -128;
       sin_table2[99] = -127;
       sin_table2[100] = -126;
       sin_table2[101] = -125;
       sin_table2[102] = -123;
       sin_table2[103] = -121;
       sin_table2[104] = -119;
       sin_table2[105] = -116;
       sin_table2[106] = -113;
       sin_table2[107] = -110;
       sin_table2[108] = -107;
       sin_table2[109] = -103;
       sin_table2[110] = -99;
       sin_table2[111] = -95;
       sin_table2[112] = -91;
       sin_table2[113] = -86;
       sin_table2[114] = -82;
       sin_table2[115] = -77;
       sin_table2[116] = -72;
       sin_table2[117] = -66;
       sin_table2[118] = -61;
       sin_table2[119] = -55;
       sin_table2[120] = -49;
       sin_table2[121] = -44;
       sin_table2[122] = -38;
       sin_table2[123] = -32;
       sin_table2[124] = -25;
       sin_table2[125] = -19;
       sin_table2[126] = -13;
       sin_table2[127] = -7;
       sin_table2[128] = -1;
       sin_table2[129] = 6;
       sin_table2[130] = 12;
       sin_table2[131] = 18;
       sin_table2[132] = 24;
       sin_table2[133] = 31;
       sin_table2[134] = 37;
       sin_table2[135] = 43;
       sin_table2[136] = 48;
       sin_table2[137] = 54;
       sin_table2[138] = 60;
       sin_table2[139] = 65;
       sin_table2[140] = 71;
       sin_table2[141] = 76;
       sin_table2[142] = 81;
       sin_table2[143] = 85;
       sin_table2[144] = 90;
       sin_table2[145] = 94;
       sin_table2[146] = 98;
       sin_table2[147] = 102;
       sin_table2[148] = 106;
       sin_table2[149] = 109;
       sin_table2[150] = 112;
       sin_table2[151] = 115;
       sin_table2[152] = 118;
       sin_table2[153] = 120;
       sin_table2[154] = 122;
       sin_table2[155] = 124;
       sin_table2[156] = 125;
       sin_table2[157] = 126;
       sin_table2[158] = 127;
       sin_table2[159] = 127;
       sin_table2[160] = 127;
       sin_table2[161] = 127;
       sin_table2[162] = 127;
       sin_table2[163] = 126;
       sin_table2[164] = 125;
       sin_table2[165] = 124;
       sin_table2[166] = 122;
       sin_table2[167] = 120;
       sin_table2[168] = 118;
       sin_table2[169] = 115;
       sin_table2[170] = 112;
       sin_table2[171] = 109;
       sin_table2[172] = 106;
       sin_table2[173] = 102;
       sin_table2[174] = 98;
       sin_table2[175] = 94;
       sin_table2[176] = 90;
       sin_table2[177] = 85;
       sin_table2[178] = 81;
       sin_table2[179] = 76;
       sin_table2[180] = 71;
       sin_table2[181] = 65;
       sin_table2[182] = 60;
       sin_table2[183] = 54;
       sin_table2[184] = 48;
       sin_table2[185] = 43;
       sin_table2[186] = 37;
       sin_table2[187] = 31;
       sin_table2[188] = 24;
       sin_table2[189] = 18;
       sin_table2[190] = 12;
       sin_table2[191] = 6;
       sin_table2[192] = 0;
       sin_table2[193] = -7;
       sin_table2[194] = -13;
       sin_table2[195] = -19;
       sin_table2[196] = -25;
       sin_table2[197] = -32;
       sin_table2[198] = -38;
       sin_table2[199] = -44;
       sin_table2[200] = -49;
       sin_table2[201] = -55;
       sin_table2[202] = -61;
       sin_table2[203] = -66;
       sin_table2[204] = -72;
       sin_table2[205] = -77;
       sin_table2[206] = -82;
       sin_table2[207] = -86;
       sin_table2[208] = -91;
       sin_table2[209] = -95;
       sin_table2[210] = -99;
       sin_table2[211] = -103;
       sin_table2[212] = -107;
       sin_table2[213] = -110;
       sin_table2[214] = -113;
       sin_table2[215] = -116;
       sin_table2[216] = -119;
       sin_table2[217] = -121;
       sin_table2[218] = -123;
       sin_table2[219] = -125;
       sin_table2[220] = -126;
       sin_table2[221] = -127;
       sin_table2[222] = -128;
       sin_table2[223] = -128;
       sin_table2[224] = -129;
       sin_table2[225] = -128;
       sin_table2[226] = -128;
       sin_table2[227] = -127;
       sin_table2[228] = -126;
       sin_table2[229] = -125;
       sin_table2[230] = -123;
       sin_table2[231] = -121;
       sin_table2[232] = -119;
       sin_table2[233] = -116;
       sin_table2[234] = -113;
       sin_table2[235] = -110;
       sin_table2[236] = -107;
       sin_table2[237] = -103;
       sin_table2[238] = -99;
       sin_table2[239] = -95;
       sin_table2[240] = -91;
       sin_table2[241] = -86;
       sin_table2[242] = -82;
       sin_table2[243] = -77;
       sin_table2[244] = -72;
       sin_table2[245] = -66;
       sin_table2[246] = -61;
       sin_table2[247] = -55;
       sin_table2[248] = -49;
       sin_table2[249] = -44;
       sin_table2[250] = -38;
       sin_table2[251] = -32;
       sin_table2[252] = -25;
       sin_table2[253] = -19;
       sin_table2[254] = -13;
       sin_table2[255] = -7;
	 end

   always @(phase) begin
	//    clk_sign           sign    
       if (phase==0)begin
		  if (correlation1 > correlation2)
           sign <= 1;
       else
           sign <= 0;
       correlation1 <= 0; // 
       correlation2 <= 0; //
		  end
		  else begin
       //    phase    signal  ı仯          
       correlation1 = correlation1 + sin_table1[phase] * signal;
       correlation2 = correlation2 + sin_table2[phase] * signal;	 
		  end 
   end

endmodule